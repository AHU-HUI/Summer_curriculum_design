/*******************************/
/***** 单个数码管译码模块 ******/
/*******************************/

// 共阳数码管
module DP1_P(
    input[3:0] num,
    output reg[6:0] data    // GFEDCBA
);

/*
    -----A-----
    |         |
    F         B
    |         |
    -----G-----
    |         |
    E         C
    |         |
    -----D-----
*/

always @(num)
case (num)
    4'b0000: data = 7'b100_0000;
    4'b0001: data = 7'b111_1001;
    4'b0010: data = 7'b010_0100;
    4'b0011: data = 7'b011_0000;
    4'b0100: data = 7'b001_1001;
    4'b0101: data = 7'b001_0010;
    4'b0110: data = 7'b000_0010;
    4'b0111: data = 7'b111_1000;
    4'b1000: data = 7'b000_0000;
    4'b1001: data = 7'b001_0000;
    4'b1010: data = 7'b000_1000;
    4'b1011: data = 7'b000_0011;
    4'b1100: data = 7'b100_0110;
    4'b1101: data = 7'b010_0001;
    4'b1110: data = 7'b000_0110;
    4'b1111: data = 7'b000_1110;
endcase

endmodule


// 共阴数码管
module DP1_N(
    input[3:0] num,
    output reg[6:0] data    // GFEDCBA
);

always @(num)
case (num)
    4'b0000: data = 7'b011_1111;
    4'b0001: data = 7'b000_0110;
    4'b0010: data = 7'b101_1011;
    4'b0011: data = 7'b100_1111;
    4'b0100: data = 7'b110_0110;
    4'b0101: data = 7'b110_1101;
    4'b0110: data = 7'b111_1101;
    4'b0111: data = 7'b000_0111;
    4'b1000: data = 7'b111_1111;
    4'b1001: data = 7'b110_1111;
    4'b1010: data = 7'b111_0111;
    4'b1011: data = 7'b111_1100;
    4'b1100: data = 7'b011_1001;
    4'b1101: data = 7'b101_1110;
    4'b1110: data = 7'b111_1001;
    4'b1111: data = 7'b111_0001;
endcase

endmodule